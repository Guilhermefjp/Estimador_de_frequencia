library verilog;
use verilog.vl_types.all;
entity exemplo1_tb is
end exemplo1_tb;
